/*
  TB file for serializer
*/

module tb_serializer ();

endmodule
