module encoder_5b6b (
  input clk,
  input reset,
  input logic [4:0] data_in,
  output logic [5:0] data_out
);

endmodule