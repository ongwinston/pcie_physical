module encoder_3b4b (
  input clk,
  input reset,
  input logic [2:0] data_in,
  output logic [3:0] data_out
);

endmodule